`timescale 1ns / 1ps

module vga_controller(
    input clk,   
    input reset,        
    output video_on,    
    output hsync,      
    output vsync,     
    output p_pixel,     
    output [9:0] x,     
    output [9:0] y     
    );
    
    // Based on VGA standards found at vesa.org for 640x480 resolution
    // Total horizontal width of screen = 800 pixels, partitioned  into sections
    parameter HD = 640;             // horizontal display area width 
    parameter HF = 48;              // horizontal front porch width 
    parameter HB = 16;              // horizontal back porch width 
    parameter HR = 96;              // horizontal retrace width 
    parameter HMAX = HD+HF+HB+HR-1; // max value of horizontal counter = 799
    // Total vertical length of screen = 525 pixels, partitioned into sections
    parameter VD = 480;             // vertical display area length 
    parameter VF = 10;              // vertical front porch length  
    parameter VB = 33;              // vertical back porch length  
    parameter VR = 2;               // vertical retrace length   
    parameter VMAX = VD+VF+VB+VR-1; // max value of vertical counter = 524   
    
	reg  [1:0] r_25MHz;
	wire w_25MHz;
	
    always @(posedge clk or posedge reset) begin
        if (reset)
            r_25MHz <= 0;
        else if (r_25MHz == 2)  // When counter reaches 2, reset it
            r_25MHz <= 0;
        else
            r_25MHz <= r_25MHz + 1;
    end

    assign w_25MHz = (r_25MHz == 2);  // w_25MHz is high when r_25MHz is 2

	
	/*always @(posedge clk or posedge reset) begin
    if (reset)
        r_25MHz <= 0;
    else if (r_25MHz == 2)  // When counter reaches 2, reset it
        r_25MHz <= 0;
    else
        r_25MHz <= r_25MHz + 1;
    end

    assign w_25MHz = (r_25MHz == 2);  // w_25MHz is high when r_25MHz is 2*/

    
    // Counter Registers, two each for buffering to avoid glitches
    reg [9:0] h_count_reg, h_count_next;
    reg [9:0] v_count_reg, v_count_next;
    
    // Output Buffers
    reg v_sync_reg, h_sync_reg;
    wire v_sync_next, h_sync_next;
    
    // Register Control
    always @(posedge clk or posedge reset)
        if(reset) begin
            v_count_reg <= 0;
            h_count_reg <= 0;
            v_sync_reg  <= 1'b0;
            h_sync_reg  <= 1'b0;
        end
        else begin
            v_count_reg <= v_count_next;
            h_count_reg <= h_count_next;
            v_sync_reg  <= v_sync_next;
            h_sync_reg  <= h_sync_next;
        end
         
   /* //Logic for horizontal counter
    always @(posedge w_25MHz or posedge reset)      // pixel tick
        if(reset)
            h_count_next = 0;
        else
            if(h_count_reg == HMAX)                 // end of horizontal scan
                h_count_next = 0;
            else
                h_count_next = h_count_reg + 1;         
  
    // Logic for vertical counter
    always @(posedge w_25MHz or posedge reset)
        if(reset)
            v_count_next = 0;
        else
            if(h_count_reg == HMAX)                 // end of horizontal scan
                if((v_count_reg == VMAX))           // end of vertical scan
                    v_count_next = 0;
                else
                    v_count_next = v_count_reg + 1;*/
        // Logic for horizontal counter
        always @(posedge w_25MHz or posedge reset) begin
            if (reset)
                h_count_next <= 0;  // Reset horizontal count
            else if (h_count_reg == HMAX)  // Check if end of horizontal scan
                h_count_next <= 0;  // Reset to zero
            else
                h_count_next <= h_count_reg + 1;  // Increment horizontal count
        end

        // Logic for vertical counter
        always @(posedge w_25MHz or posedge reset) begin
            if (reset)
                v_count_next <= 0;  // Reset vertical count
            else if (h_count_reg == HMAX) begin
                if (v_count_reg == VMAX)  // Check if end of vertical scan
                    v_count_next <= 0;  // Reset to zero
                else
                    v_count_next <= v_count_reg + 1;  // Increment vertical count
            end
        end



        
    // h_sync_next asserted within the horizontal retrace area
    assign h_sync_next = (h_count_reg >= (HD+HB) && h_count_reg <= (HD+HB+HR-1));
    
    // v_sync_next asserted within the vertical retrace area
    assign v_sync_next = (v_count_reg >= (VD+VB) && v_count_reg <= (VD+VB+VR-1));
    
    // Video ON/OFF - only ON while pixel counts are within the display area
    assign video_on = (h_count_reg < HD) && (v_count_reg < VD); // 0-639 and 0-479 
            
    // Outputs
    assign hsync  = h_sync_reg;
    assign vsync  = v_sync_reg;
    assign x      = h_count_reg;
    assign y      = v_count_reg;
    assign p_pixel = w_25MHz;
            
endmodule
